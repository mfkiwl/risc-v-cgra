
`include "LocalBus.v"
`timescale 1ns / 1ps

module tb_local_bus_top;

    // Inputs to the local_bus_top module
    reg clk;
    reg reset;
    reg [31:0] global_mem_read_data; // Data read from global memory
    reg global_mem_ack;             // Acknowledgment signal from global memory

    // Outputs from the local_bus_top module
    wire [31:0] global_mem_address;       // Address for global memory operations
    wire [31:0] global_mem_write_data;    // Data to write to global memory
    wire global_mem_write;                // Write enable signal for global memory
    wire global_mem_read;                 // Read enable signal for global memory
    wire [127:0] result_out;              // Result output from the cluster

    // Instantiate the local_bus_top module
    local_bus_top uut (
        .clk(clk),
        .reset(reset),
        .global_mem_address(global_mem_address),
        .global_mem_write_data(global_mem_write_data),
        .global_mem_read_data(global_mem_read_data),
        .global_mem_ack(global_mem_ack),
        .global_mem_write(global_mem_write),
        .global_mem_read(global_mem_read),
        .result_out(result_out)
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // Clock period = 10 time units
    end

    // Testbench logic
    initial begin
        // Dump waveform for debugging
        $dumpfile("tb_local_bus_top.vcd");
        $dumpvars(0, tb_local_bus_top);

        // Initialize input signals
        reset = 1;
        global_mem_read_data = 32'b0;
        global_mem_ack = 0;

        #10 reset = 0; // Release reset

        //Need time to load instructions and wait for responses from PEs

        // Test Case 1: Initialize global memory read operation
        $display("Test Case 1: Global memory read operation");
        global_mem_ack = 1;
        #10 global_mem_ack = 0;

        // Test Case 2: Global memory write operation
        $display("Test Case 2: Global memory write operation");
        global_mem_read_data = 32'hCAFEBABE; // Mock data from global memory
        global_mem_ack = 1; // Acknowledge global memory
        #10 global_mem_ack = 0;

        // Test Case 3: Simulate PE requests and grant arbitration
        $display("Test Case 3: Simulate PE bus requests and arbitration");
        // Simulate requests from the PEs and check grant signals
        // For example:
        // bus_request signals will be generated by the PE interfaces
        // Ensure the arbiter properly handles grant signal assignments

        #50;

        // Test Case 4: Reset the cluster
        $display("Test Case 4: Reset cluster components");
        reset = 1;
        #10 reset = 0;

        // End simulation
        $finish;
    end

endmodule
